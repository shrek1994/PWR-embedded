library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

package utills is
    type data_type is array (0 to 31) of std_logic_vector (8 downto 0);
end package utills;

package body utills is

end utills;
